module xor_1 (A,B,O);
	input A;
	input B;
	output C;
	xor G1(O,A,B);
endmodule


