library verilog;
use verilog.vl_types.all;
entity Sin_t_tb is
end Sin_t_tb;
