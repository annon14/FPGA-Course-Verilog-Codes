`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:54:27 04/19/2017 
// Design Name: 
// Module Name:    Top_module 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Top_module( 
    );
	Shift_reg_8bit ins1 () ;
	shift_reg_8bit #12 ins1();
	shift_reg_8bit #12 ins1();
	shift_reg_8bit ins1.w = 12 ;
	

endmodule
