`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:48:28 03/08/2017 
// Design Name: 
// Module Name:    full_adder_8bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module full_adder( A , B , Cin , Cout ,Sum )
    );
 input  A ;
 input  B ;
 input Cin ;
 output Sum ; 
 output Cout ;
    
endmodule
